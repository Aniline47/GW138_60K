`define module_name DDS_II_DA
